module btb #(
    parameter SETS = 8,
    parameter WAYS = 2,
    parameter TAGW = 27
)(
    input              clk,
    input              rst,

    // ================= FETCH =================
    input      [31:0]  pc,
    output reg         predict_valid,
    output reg         predict_taken,
    output reg [31:0]  predict_target,

    // ================= UPDATE =================
    input              update_en,
    input      [29:0]  update_pc,
    input              actual_taken,
    input      [31:0]  update_target
);

    // ============================================================
    // FETCH STAGE
    // ============================================================
    wire [2:0] fetch_set; // WHAT: BTB set index WHY: Selects one set in 2-way BTB HOW: Derived from PC bits WHEN: BTB lookup
 //   wire [TAGW-1:0] fetch_tag;
    wire hit0, hit1; // WHAT: Way hit signals WHY: Identify matching BTB entry HOW: Tag compare logic WHEN: Fetch lookup

    // Data returned from btb_file for fetch read
    wire rd_valid0, rd_valid1; // WHAT: Valid bits for each way WHY: Ignore empty entries HOW: Stored in BTB file WHEN: Read stage
    wire [TAGW-1:0] rd_tag0, rd_tag1; // WHAT: Stored tags WHY: Used for tag comparison HOW: Read from BTB arrays WHEN: Fetch lookup
    wire [31:0] rd_target0, rd_target1; // WHAT: Stored branch targets WHY: Used for predicted PC HOW: Read from BTB WHEN: BTB hit
    wire [1:0]  rd_state0, rd_state1; // WHAT: 2-bit predictor states WHY: Predict taken/not-taken HOW: Saturating counter bits WHEN: Prediction
    wire rd_lru; // WHAT: LRU bit for set WHY: Select replacement way HOW: Stored per set WHEN: On BTB update

    // ----------------- FETCH READ MODULE -----------------
    btb_read #(.TAGW(TAGW)) U_READ (
        .pc(pc[31:2]),

        .rd_valid0(rd_valid0),
        .rd_tag0(rd_tag0),

        .rd_valid1(rd_valid1),
        .rd_tag1(rd_tag1),

        .set_index(fetch_set),
      //  .tag(fetch_tag),
        .hit0(hit0),
        .hit1(hit1)
    );

    // ----------------- FETCH OUTPUT LOGIC -----------------
    always @(hit0 or hit1 or rd_state0[1] or  rd_state1[1] or rd_target0 or rd_target1 or pc) begin
        predict_valid = hit0 | hit1; // WHAT: Indicate BTB hit WHY: Enable use of prediction HOW: OR of both way hits WHEN: Fetch stage

        if (hit0) begin
            predict_taken  = rd_state0[1]; // WHAT: Predicted direction from way0 WHY: Use MSB of state HOW: State bit check WHEN: Way0 hit
            predict_target = rd_target0; // WHAT: Predicted target from way0 WHY: Jump to correct address HOW: Read target mux WHEN: Way0 hit
        end
        else if (hit1) begin
            predict_taken  = rd_state1[1]; // WHAT: Predicted direction from way1 WHY: Use MSB of state HOW: State bit check WHEN: Way1 hit
            predict_target = rd_target1; // WHAT: Predicted target from way1 WHY: Jump to correct address HOW: Read target mux WHEN: Way1 hit
        end
        else begin
            predict_taken  = 1'b0; // WHAT: Default not-taken prediction WHY: No BTB entry found HOW: Force zero WHEN: BTB miss
            predict_target = pc + 32'd4; // WHAT: Sequential target WHY: Continue normal flow HOW: PC+4 WHEN: No prediction
        end
    end

    // ============================================================
    // UPDATE STAGE (WRITE PATH)
    // ============================================================
   // wire [2:0] upd_set = update_pc[2:0];
   // wire [TAGW-1:0] upd_tag = update_pc[29:3];

    // Signals from BTB file for update side read
    wire upd_valid0 = rd_valid0; // WHAT: Valid bit of way0 for update WHY: Check if entry exists HOW: Reuse fetch read data WHEN: Update stage
    wire upd_valid1 = rd_valid1; // WHAT: Valid bit of way1 for update WHY: Check if entry exists HOW: Reuse fetch read data WHEN: Update stage
    wire [TAGW-1:0] upd_tag0 = rd_tag0; // WHAT: Tag of way0 for update WHY: Match update PC HOW: Reuse tag read WHEN: Update stage
    wire [TAGW-1:0] upd_tag1 = rd_tag1; // WHAT: Tag of way1 for update WHY: Match update PC HOW: Reuse tag read WHEN: Update stage

    // Predictor states for write logic
  //  wire [1:0] next_state0, next_state1;

    // ----------------- WRITE CONTROL -----------------
    wire         wr_en; // WHAT: Write enable for BTB file WHY: Control update operation HOW: Generated by update logic WHEN: Branch resolved
    wire [2:0]   wr_set; // WHAT: Set index to write WHY: Select correct BTB set HOW: From update PC bits WHEN: BTB update
    wire         wr_way; // WHAT: Selected way to write WHY: Choose hit or replacement way HOW: LRU or hit select WHEN: Update stage
    wire         wr_valid; // WHAT: Valid bit to write WHY: Mark entry as valid HOW: Set to 1 on allocation WHEN: New entry
    wire [TAGW-1:0] wr_tag; // WHAT: Tag to write WHY: Identify branch PC HOW: From update PC WHEN: BTB update
    wire [31:0] wr_target; // WHAT: Target address to write WHY: Future prediction target HOW: From resolved jump WHEN: Branch taken
    wire [1:0]  wr_state; // WHAT: New predictor state WHY: Update branch history HOW: FSM update logic WHEN: After branch resolution

    wire wr_lru_en; // WHAT: LRU update enable WHY: Maintain replacement policy HOW: Set on BTB access/update WHEN: After update
    wire wr_lru_val; // WHAT: New LRU value WHY: Mark recently used way HOW: Write to LRU bit WHEN: Update stage

    // ----------------- UPDATE MODULE -----------------
    btb_write #(.TAGW(TAGW)) U_WRITE (
        .clk(clk),
        .rst(rst),
        .update_en(update_en),
        .update_pc(update_pc),
        .actual_taken(actual_taken),
        .update_target(update_target),

        .rd_valid0_upd(upd_valid0),
        .rd_tag0_upd(upd_tag0),
        .rd_valid1_upd(upd_valid1),
        .rd_tag1_upd(upd_tag1),
        .rd_lru_upd(rd_lru),

        .wr_en(wr_en),
        .wr_set(wr_set),
        .wr_way(wr_way),
        .wr_valid(wr_valid),
        .wr_tag(wr_tag),
        .wr_target(wr_target),
        .wr_state(wr_state),

        .wr_lru_en(wr_lru_en),
        .wr_lru_val(wr_lru_val),

        .state0_in(rd_state0),
        .state1_in(rd_state1)
     //  .next_state0(next_state0),
     //  .next_state1(next_state1)
    );

    // ============================================================
    // BTB FILE (Storage Arrays)
    // ============================================================

    btb_file #(.SETS(SETS), .WAYS(WAYS), .TAGW(TAGW)) U_FILE (
        .clk(clk),
        .rst(rst),

        // READ side
        .rd_set(fetch_set),
      //  .rd_way0(1'b0),
        .rd_valid0(rd_valid0),
        .rd_tag0(rd_tag0),
        .rd_target0(rd_target0),
        .rd_state0(rd_state0),

    //    .rd_way1(1'b0),
        .rd_valid1(rd_valid1),
        .rd_tag1(rd_tag1),
        .rd_target1(rd_target1),
        .rd_state1(rd_state1),

        .rd_lru(rd_lru),

        // WRITE side
        .wr_en(wr_en),
        .wr_set(wr_set),
        .wr_way(wr_way),
        .wr_valid(wr_valid),
        .wr_tag(wr_tag),
        .wr_target(wr_target),
        .wr_state(wr_state),

        .wr_lru_en(wr_lru_en),
        .wr_lru_val(wr_lru_val)
    );

endmodule

